   ,max_ep ,max_it ,batch ,datas ,LR    ,ue  ,train_t ,res_waste ,rew    ,pred_tt ,er_prc_tt ,er_abs_tt ,pred_rew ,er_prc_rew ,er_abs_rew ,pred_rw ,er_prc_rw ,er_abs_rw
12 ,     1 ,     2 ,  123 ,22349 ,0.031 ,  5 , 10.314 ,  905.618 ,-2.007 ,  1.996 ,   80.5   ,-8.317    ,-3.164   ,    58.25  ,-1.157     ,357.537 ,   60.5   ,-548.081
 0 ,     1 ,     2 ,   21 ,19761 ,0.007 ,  3 , 10.098 ,  883.486 ,-2.014 ,  2.568 ,   74.5   ,-7.531    ,-2.282   ,    14.0   ,-0.268     ,142.555 ,   83.75  ,-740.931
 3 ,     1 ,     2 ,   99 ,22953 ,0.028 , 98 , 10.036 ,  891.777 ,-2.004 ,  1.634 ,   83.75  ,-8.402    ,-4.019   ,   102.25  ,-2.015     ,507.689 ,   43.25  ,-384.088
14 ,     1 ,     2 ,  129 ,22612 ,0.009 ,  4 ,  9.964 ,  917.789 ,-1.945 ,  2.101 ,   79.0   ,-7.864    ,-2.878   ,    48.25  ,-0.933     ,314.346 ,   65.75  ,-603.443
 5 ,     1 ,     2 ,  103 ,22593 ,0.109 ,  3 ,  9.896 ,  903.942 ,-1.961 ,  1.646 ,   83.25  ,-8.25     ,-3.791   ,    96.25  ,-1.83      ,503.889 ,   44.0   ,-400.053
29 ,     1 ,     2 ,  204 ,25383 ,0.011 ,  1 ,  9.838 ,  891.522 ,-1.882 ,  1.092 ,   89.0   ,-8.746    ,-2.375   ,    27.25  ,-0.493     ,742.998 ,   16.5   ,-148.524
24 ,     1 ,     2 ,  186 ,20542 ,0.001 ,  3 ,  9.79  ,  896.191 ,-1.962 ,  1.431 ,   85.25  ,-8.359    ,-2.392   ,    22.75  ,-0.43      ,601.13  ,   33.0   ,-295.06
11 ,     1 ,     2 ,  120 ,19795 ,0.003 ,  9 ,  9.712 ,  924.471 ,-1.887 ,  1.945 ,   79.75  ,-7.767    ,-3.283   ,    74.0   ,-1.396     ,386.644 ,   58.25  ,-537.827
37 ,    77 ,     2 ,  100 ,20352 ,0.006 ,  5 ,  9.661 ,  917.022 ,-2.252 ,  1.599 ,   82.794 ,-8.062    ,-3.681   ,    96.676 ,-1.429     ,530.394 ,   41.941 ,-386.628
13 ,     1 ,     2 ,  129 ,22599 ,0.059 ,  1 ,  9.616 ,  871.879 ,-1.924 ,  2.101 ,   78.0   ,-7.515    ,-2.977   ,    55.0   ,-1.053     ,317.082 ,   63.75  ,-554.796
 2 ,     1 ,     2 ,   30 ,23158 ,0.006 , 66 ,  9.413 ,  874.85  ,-1.759 ,  2.468 ,   73.75  ,-6.945    ,-2.102   ,    20.0   ,-0.343     ,150.671 ,   83.0   ,-724.179
 7 ,     1 ,     2 ,  107 ,23236 ,0.006 ,  5 ,  9.403 ,  937.783 ,-1.836 ,  1.716 ,   81.25  ,-7.687    ,-3.518   ,    96.0   ,-1.681     ,473.562 ,   49.75  ,-464.221
16 ,     1 ,     2 ,  138 ,18587 ,0.001 , 46 ,  9.391 ,  888.164 ,-1.741 ,  2.261 ,   76.0   ,-7.13     ,-2.632   ,    51.5   ,-0.89      ,254.533 ,   71.25  ,-633.631
28 ,     1 ,     2 ,  195 ,19816 ,0.029 ,  4 ,  9.341 ,  894.866 ,-1.796 ,  1.173 ,   87.75  ,-8.168    ,-2.468   ,    38.25  ,-0.672     ,706.6   ,   21.0   ,-188.266
27 ,     1 ,     2 ,  194 ,23379 ,0.013 , 57 ,  9.284 ,  874.984 ,-1.797 ,  1.199 ,   87.0   ,-8.085    ,-2.431   ,    36.0   ,-0.634     ,697.187 ,   20.25  ,-177.796
15 ,     1 ,     2 ,  133 ,23285 ,0.028 , 87 ,  9.228 ,  895.427 ,-1.776 ,  2.172 ,   76.5   ,-7.056    ,-3.007   ,    70.75  ,-1.231     ,286.026 ,   68.25  ,-609.401
34 ,    30 ,     2 ,   23 ,25380 ,0.008 ,  3 ,  9.171 ,  912.491 ,-2.144 ,  2.538 ,   71.25  ,-6.633    ,-2.393   ,    59.2   ,-0.248     ,140.373 ,   84.55  ,-772.119
 4 ,     1 ,     2 ,  100 ,22605 ,0.003 , 66 ,  9.165 ,  920.916 ,-1.791 ,  1.592 ,   82.25  ,-7.572    ,-3.995   ,   124.75  ,-2.204     ,529.732 ,   42.0   ,-391.184
 1 ,     1 ,     2 ,   30 ,22559 ,0.01  ,  3 ,  9.149 ,  893.064 ,-1.815 ,  2.469 ,   71.75  ,-6.68     ,-2.078   ,    36.25  ,-0.263     ,148.149 ,   83.25  ,-744.914
19 ,     1 ,     2 ,  153 ,22935 ,0.017 ,  5 ,  9.093 ,  910.547 ,-1.716 ,  2.381 ,   73.75  ,-6.712    ,-2.24    ,    32.0   ,-0.524     ,203.531 ,   77.75  ,-707.016
35 ,    30 ,     2 ,  114 ,19771 ,0.027 , 16 ,  9.086 ,  915.181 ,-2.088 ,  1.844 ,   78.738 ,-7.242    ,-3.441   ,   132.357 ,-1.353     ,419.224 ,   54.0   ,-495.957
 6 ,     1 ,     2 ,  105 ,21294 ,0.009 , 14 ,  9.072 ,  891.892 ,-1.856 ,  1.683 ,   81.25  ,-7.39     ,-3.618   ,    96.0   ,-1.762     ,486.219 ,   45.5   ,-405.673
18 ,     1 ,     2 ,  152 ,20470 ,0.013 , 49 ,  9.069 ,  892.754 ,-1.798 ,  2.412 ,   73.0   ,-6.658    ,-2.209   ,    26.75  ,-0.41      ,190.312 ,   78.75  ,-702.441
23 ,     1 ,     2 ,  185 ,21707 ,0.003 , 14 ,  8.994 ,  920.158 ,-1.76  ,  1.458 ,   83.25  ,-7.535    ,-2.512   ,    56.0   ,-0.752     ,591.333 ,   35.75  ,-328.826
26 ,     1 ,     2 ,  192 ,19783 ,0.032 , 14 ,  8.953 ,  930.614 ,-1.709 ,  1.26  ,   85.75  ,-7.693    ,-2.494   ,    50.75  ,-0.785     ,669.681 ,   28.0   ,-260.933
33 ,    10 ,     2 ,  111 ,22355 ,0.029 ,  1 ,  8.894 ,  934.595 ,-2.0   ,  1.788 ,   79.05  ,-7.106    ,-3.594   ,   138.375 ,-1.593     ,440.966 ,   52.475 ,-493.629
 8 ,     1 ,     2 ,  110 ,22602 ,0.017 , 44 ,  8.873 ,  916.783 ,-1.738 ,  1.768 ,   80.25  ,-7.105    ,-3.559   ,   105.75  ,-1.821     ,453.36  ,   50.5   ,-463.422
30 ,     1 ,     2 ,  205 ,19794 ,0.003 , 55 ,  8.861 ,  959.783 ,-1.706 ,  1.105 ,   87.5   ,-7.756    ,-2.52    ,    49.75  ,-0.814     ,743.737 ,   22.25  ,-216.046
 9 ,     1 ,     2 ,  114 ,25403 ,0.011 ,  5 ,  8.848 ,  907.949 ,-1.739 ,  1.842 ,   78.5   ,-7.006    ,-3.252   ,    92.0   ,-1.513     ,425.314 ,   53.0   ,-482.635
22 ,     1 ,     2 ,  182 ,23226 ,0.003 ,100 ,  8.783 ,  927.047 ,-1.757 ,  1.544 ,   82.0   ,-7.238    ,-2.66    ,    52.75  ,-0.903     ,556.307 ,   40.0   ,-370.741
17 ,     1 ,     2 ,  139 ,22428 ,0.029 , 80 ,  8.635 ,  896.982 ,-1.503 ,  2.276 ,   73.0   ,-6.358    ,-2.811   ,   107.0   ,-1.308     ,242.719 ,   73.0   ,-654.263
10 ,     1 ,     2 ,  118 ,22600 ,0.154 ,  2 ,  8.633 ,  896.785 ,-1.6   ,  1.908 ,   77.25  ,-6.725    ,-3.327   ,   131.0   ,-1.726     ,395.949 ,   55.75  ,-500.836
25 ,     1 ,     2 ,  189 ,19777 ,0.031 ,  1 ,  8.251 ,  935.688 ,-1.553 ,  1.347 ,   83.0   ,-6.905    ,-2.476   ,    69.25  ,-0.922     ,632.735 ,   32.25  ,-302.953
36 ,    30 ,     2 ,  191 ,20290 ,0.005 , 48 ,  8.244 ,  927.978 ,-1.744 ,  1.289 ,   83.622 ,-6.956    ,-2.341   ,   229.622 ,-0.596     ,657.776 ,   28.778 ,-270.202
20 ,     1 ,     2 ,  155 ,20069 ,0.008 , 14 ,  8.232 ,  912.693 ,-1.627 ,  2.327 ,   71.25  ,-5.905    ,-2.218   ,    40.0   ,-0.59      ,223.665 ,   75.25  ,-689.028
31 ,     1 ,     2 ,  232 ,25403 ,0.006 , 13 ,  8.034 ,  911.941 ,-1.426 ,  1.53  ,   80.25  ,-6.504    ,-2.346   ,    86.0   ,-0.92      ,568.253 ,   37.5   ,-343.688
21 ,     1 ,     2 ,  167 ,20058 ,0.022 ,  1 ,  7.936 ,  936.555 ,-1.631 ,  1.98  ,   74.75  ,-5.956    ,-2.33    ,    44.0   ,-0.699     ,370.907 ,   60.25  ,-565.648
32 ,     1 ,     2 ,  273 ,23415 ,0.129 ,  7 ,  7.758 ,  920.227 ,-1.332 ,  2.166 ,   71.5   ,-5.592    ,-2.366   ,    99.0   ,-1.034     ,314.439 ,   65.75  ,-605.788
