,max_ep,max_it,batch,datas,LR,ue,train_t,res_waste,rew,pred_tt,er_prc_tt,er_abs_tt,pred_rew,er_prc_rew,er_abs_rew,pred_rw,er_prc_rw,er_abs_rw
0,100,5,100,50000,0.01,10,5.769,659.326,-1.993,4.454,21.373,-1.316,-3.888,150.294,-1.896,733.906,12.542,74.579
