   ,max_ep ,max_it ,batch ,datas ,LR    ,ue  ,train_t ,res_waste ,rew    ,pred_tt ,er_prc_tt ,er_abs_tt ,pred_rew ,er_prc_rew ,er_abs_rew ,pred_rw ,er_prc_rw ,er_abs_rw
 1 ,     1 ,     1 ,   30 ,22698 ,0.005 ,  5 ,  2.081 ,  115.257 ,-1.608 ,  2.925 ,   40.5   ,0.843     ,-1.796   ,    45.25  ,-0.189     ,160.144 ,   39.0   ,44.887
28 ,     2 ,     1 ,   30 , 4226 ,0.005 ,  5 ,  2.107 ,  111.552 ,-2.002 ,  2.934 ,   39.25  ,0.827     ,-1.753   ,    24.625 ,0.249      ,195.668 ,   75.75  ,84.115
 2 ,     1 ,     1 ,   30 ,23756 ,0.005 ,  5 ,  2.118 ,  111.263 ,-1.827 ,  2.926 ,   38.25  ,0.807     ,-1.771   ,    24.75  ,0.056      ,159.792 ,   44.0   ,48.53
36 ,     8 ,     1 ,   30 ,20725 ,0.005 ,  5 ,  2.146 ,  117.845 ,-2.184 ,  2.935 ,   36.906 ,0.789     ,-1.732   ,    31.969 ,0.452      ,195.062 ,   66.062 ,77.218
 0 ,     1 ,     1 ,   30 , 1898 ,0.005 ,  5 ,  2.159 ,  113.794 ,-1.598 ,  2.927 ,   35.5   ,0.768     ,-1.797   ,    19.75  ,-0.199     ,160.015 ,   40.75  ,46.221
45 ,    30 ,     1 ,   30 ,25151 ,0.005 ,  5 ,  2.164 ,  121.459 ,-2.21  ,  2.929 ,   35.81  ,0.765     ,-1.726   ,    95.143 ,0.485      ,158.176 ,   31.143 ,36.718
43 ,    30 ,     1 ,   30 ,17882 ,0.005 ,  5 ,  2.185 ,  122.551 ,-2.129 ,  2.929 ,   34.375 ,0.744     ,-1.735   ,    30.525 ,0.395      ,158.273 ,   31.025 ,35.722
38 ,    16 ,     1 ,   30 , 4759 ,0.005 ,  5 ,  2.189 ,  120.704 ,-2.263 ,  2.937 ,   34.512 ,0.747     ,-1.723   ,    33.073 ,0.54       ,196.348 ,   63.927 ,75.644
42 ,    30 ,     1 ,   30 , 1000 ,0.005 ,  5 ,  2.19  ,  120.623 ,-2.232 ,  2.898 ,   32.725 ,0.708     ,-1.915   ,    22.525 ,0.317      ,162.755 ,   36.15  ,42.132
39 ,    24 ,     1 ,   30 , 2575 ,0.005 ,  5 ,  2.19  ,  121.375 ,-2.228 ,  2.937 ,   34.575 ,0.747     ,-1.727   ,    29.7   ,0.501      ,196.386 ,   63.675 ,75.011
44 ,    30 ,     1 ,   30 ,19478 ,0.005 ,  5 ,  2.193 ,  123.026 ,-2.221 ,  2.93  ,   33.95  ,0.737     ,-1.724   ,    33.375 ,0.497      ,158.314 ,   30.05  ,35.289
40 ,    28 ,     1 ,   30 , 3383 ,0.005 ,  5 ,  2.198 ,  126.133 ,-2.296 ,  2.936 ,   33.85  ,0.738     ,-1.719   ,    32.575 ,0.577      ,194.473 ,   55.875 ,68.34
31 ,     4 ,     1 ,   30 ,25052 ,0.005 ,  5 ,  2.566 ,  186.079 ,-1.622 ,  2.947 ,   15.125 ,0.381     ,-1.795   ,    35.875 ,-0.173     ,200.021 ,    7.438 ,13.942
30 ,     4 ,     1 ,   30 , 2656 ,0.005 ,  5 ,  2.588 ,  190.582 ,-1.69  ,  2.948 ,   14.188 ,0.36      ,-1.787   ,    35.562 ,-0.098     ,200.417 ,    5.625 ,9.836
32 ,     5 ,     1 ,   30 ,23879 ,0.005 ,  5 ,  2.612 ,  188.71  ,-1.819 ,  2.946 ,   13.35  ,0.335     ,-1.768   ,    50.9   ,0.051      ,179.302 ,    4.9   ,-9.408
35 ,     8 ,     1 ,   30 ,16991 ,0.005 ,  5 ,  2.652 ,  190.772 ,-1.867 ,  2.95  ,   12.0   ,0.298     ,-1.768   ,    31.094 ,0.099      ,201.481 ,    5.875 ,10.709
53 ,    42 ,     1 ,   30 , 4007 ,0.005 ,  5 ,  2.708 ,  193.878 ,-1.969 ,  2.951 ,    9.628 ,0.243     ,-1.756   ,    39.86  ,0.213      ,200.537 ,    7.953 ,6.659
41 ,    28 ,     2 ,   30 , 3031 ,0.005 ,  5 ,  3.135 ,  261.777 ,-2.024 ,  3.549 ,   14.409 ,0.414     ,-1.675   ,    48.614 ,0.349      ,224.182 ,   14.023 ,-37.595
33 ,     6 ,     2 ,   30 , 4786 ,0.005 ,  5 ,  3.143 ,  260.034 ,-2.093 ,  3.549 ,   14.731 ,0.406     ,-1.667   ,    38.385 ,0.426      ,222.096 ,   14.5   ,-37.938
34 ,     7 ,     2 ,   30 , 1099 ,0.005 ,  5 ,  3.152 ,  264.697 ,-2.045 ,  3.549 ,   14.4   ,0.398     ,-1.673   ,    47.733 ,0.372      ,222.363 ,   15.8   ,-42.335
47 ,    30 ,     2 ,   30 , 1885 ,0.005 ,  5 ,  3.153 ,  263.317 ,-2.031 ,  3.544 ,   13.674 ,0.39      ,-1.671   ,    40.279 ,0.36       ,188.433 ,   28.279 ,-74.884
 6 ,     1 ,     2 ,   30 , 1296 ,0.005 ,  5 ,  3.263 ,  292.397 ,-1.66  ,  3.514 ,   58.8   ,0.251     ,-1.709   ,    21.4   ,-0.049     ,178.979 ,   50.4   ,-113.419
 5 ,     1 ,     2 ,   29 , 1000 ,0.005 ,  5 ,  3.492 ,  285.678 ,-1.577 ,  3.456 ,   63.0   ,-0.036    ,-2.598   ,    74.0   ,-1.021     ,172.285 ,   51.0   ,-113.393
29 ,     2 ,     2 ,   30 , 1913 ,0.005 ,  5 ,  3.563 ,  286.576 ,-2.184 ,  3.522 ,   61.9   ,-0.041    ,-1.66    ,    23.7   ,0.524      ,214.333 ,   76.4   ,-72.243
46 ,    30 ,     2 ,   30 , 1001 ,0.004 ,  5 ,  3.57  ,  303.054 ,-2.085 ,  3.515 ,   57.824 ,-0.055    ,-1.901   ,    37.588 ,0.184      ,184.273 ,   50.784 ,-118.781
48 ,    30 ,     2 ,   30 , 4567 ,0.005 ,  5 ,  3.694 ,  282.428 ,-2.008 ,  3.516 ,   59.04  ,-0.178    ,-1.681   ,    44.38  ,0.328      ,176.575 ,   46.84  ,-105.853
 7 ,     1 ,     2 ,   30 , 3255 ,0.005 ,  5 ,  3.698 ,  286.025 ,-1.544 ,  3.514 ,   60.2   ,-0.184    ,-1.741   ,    29.4   ,-0.196     ,178.531 ,   53.0   ,-107.493
 3 ,     1 ,     2 ,    1 , 1000 ,0.005 ,  5 ,  3.9   ,  275.61  ,-1.786 ,  3.602 ,   65.8   ,-0.297    ,-2.132   ,    21.8   ,-0.346     ,175.173 ,   48.6   ,-100.436
52 ,    40 ,     1 ,  150 ,24026 ,0.005 ,  5 ,  4.62  ,  375.987 ,-1.888 ,  3.012 ,   32.82  ,-1.609    ,-1.955   ,   101.12  ,-0.067     ,207.948 ,   44.5   ,-168.039
51 ,    39 ,     2 ,  150 , 1566 ,0.005 ,  5 ,  6.582 ,  620.745 ,-1.889 ,  3.652 ,   42.278 ,-2.93     ,-1.883   ,    62.204 ,0.007      ,255.328 ,   58.537 ,-365.417
27 ,     1 ,     2 ,  232 ,25403 ,0.006 , 13 ,  8.034 ,  911.941 ,-1.426 ,  2.928 ,   61.75  ,-5.106    ,-2.985   ,   137.0   ,-1.559     ,480.394 ,   47.25  ,-431.547
50 ,    30 ,     2 ,  191 ,20290 ,0.005 , 48 ,  8.244 ,  927.978 ,-1.744 ,  2.896 ,   63.178 ,-5.348    ,-2.149   ,   209.333 ,-0.405     ,482.37  ,   47.778 ,-445.608
21 ,     1 ,     2 ,  189 ,19777 ,0.031 ,  1 ,  8.251 ,  935.688 ,-1.553 ,  2.896 ,   64.0   ,-5.355    ,-2.732   ,    86.5   ,-1.179     ,488.517 ,   47.75  ,-447.17
54 ,    77 ,     2 ,  100 ,20352 ,0.006 ,  5 ,  8.571 ,  985.475 ,-1.918 ,  2.858 ,   66.25  ,-5.712    ,-3.743   ,   108.0   ,-1.826     ,633.61  ,   35.25  ,-351.864
16 ,     1 ,     2 ,  139 ,22428 ,0.029 , 80 ,  8.635 ,  896.982 ,-1.503 ,  2.858 ,   66.25  ,-5.777    ,-2.825   ,   107.75  ,-1.322     ,474.54  ,   47.0   ,-422.442
18 ,     1 ,     2 ,  182 ,23226 ,0.003 ,100 ,  8.783 ,  927.047 ,-1.757 ,  2.844 ,   67.0   ,-5.939    ,-2.526   ,    45.0   ,-0.769     ,486.866 ,   47.5   ,-440.181
26 ,     1 ,     2 ,  205 ,19794 ,0.003 , 55 ,  8.861 ,  959.783 ,-1.706 ,  2.836 ,   67.5   ,-6.025    ,-2.405   ,    43.0   ,-0.7       ,499.444 ,   47.75  ,-460.339
37 ,    10 ,     2 ,  111 ,22355 ,0.029 ,  1 ,  8.894 ,  934.595 ,-2.0   ,  2.835 ,   66.775 ,-6.059    ,-1.941   ,    56.15  ,0.059      ,487.037 ,   47.575 ,-447.558
22 ,     1 ,     2 ,  192 ,19783 ,0.032 , 14 ,  8.953 ,  930.614 ,-1.709 ,  2.827 ,   68.0   ,-6.126    ,-2.384   ,    44.25  ,-0.676     ,487.821 ,   47.5   ,-442.793
19 ,     1 ,     2 ,  185 ,21707 ,0.003 , 14 ,  8.994 ,  920.158 ,-1.76  ,  2.823 ,   67.5   ,-6.171    ,-2.303   ,    43.5   ,-0.543     ,483.702 ,   47.5   ,-436.456
49 ,    30 ,     2 ,  114 ,19771 ,0.027 , 16 ,  9.086 ,  915.181 ,-2.088 ,  2.818 ,   67.619 ,-6.267    ,-1.771   ,    58.286 ,0.317      ,479.147 ,   47.476 ,-436.034
17 ,     1 ,     2 ,  153 ,22935 ,0.017 ,  5 ,  9.093 ,  910.547 ,-1.716 ,  2.814 ,   69.0   ,-6.28     ,-2.372   ,    39.5   ,-0.656     ,480.922 ,   47.0   ,-429.625
10 ,     1 ,     2 ,  100 ,22605 ,0.003 , 66 ,  9.165 ,  920.916 ,-1.791 ,  2.845 ,   69.0   ,-6.32     ,-3.736   ,   110.5   ,-1.946     ,621.679 ,   32.25  ,-299.237
15 ,     1 ,     2 ,  133 ,23285 ,0.028 , 87 ,  9.228 ,  895.427 ,-1.776 ,  2.801 ,   69.5   ,-6.427    ,-2.289   ,    29.75  ,-0.513     ,474.165 ,   47.25  ,-421.262
23 ,     1 ,     2 ,  194 ,23379 ,0.013 , 57 ,  9.284 ,  874.984 ,-1.797 ,  2.795 ,   69.75  ,-6.488    ,-2.232   ,    25.0   ,-0.436     ,466.121 ,   47.0   ,-408.863
24 ,     1 ,     2 ,  195 ,19816 ,0.029 ,  4 ,  9.341 ,  894.866 ,-1.796 ,  2.79  ,   70.0   ,-6.552    ,-2.251   ,    26.0   ,-0.454     ,473.732 ,   47.0   ,-421.134
11 ,     1 ,     2 ,  107 ,23236 ,0.006 ,  5 ,  9.403 ,  937.783 ,-1.836 ,  2.784 ,   69.75  ,-6.619    ,-2.217   ,    23.5   ,-0.38      ,491.646 ,   47.75  ,-446.137
 8 ,     1 ,     2 ,   30 ,23158 ,0.006 , 66 ,  9.413 ,  874.85  ,-1.759 ,  3.727 ,   60.5   ,-5.686    ,-1.938   ,    10.5   ,-0.179     ,245.883 ,   71.75  ,-628.967
12 ,     1 ,     2 ,  120 ,19795 ,0.003 ,  9 ,  9.712 ,  924.471 ,-1.887 ,  2.754 ,   71.75  ,-6.958    ,-2.056   ,     9.0   ,-0.169     ,485.431 ,   47.5   ,-439.04
20 ,     1 ,     2 ,  186 ,20542 ,0.001 ,  3 ,  9.79  ,  896.191 ,-1.962 ,  2.746 ,   71.5   ,-7.044    ,-1.873   ,     6.75  ,0.088      ,474.543 ,   47.0   ,-421.648
25 ,     1 ,     2 ,  204 ,25383 ,0.011 ,  1 ,  9.838 ,  891.522 ,-1.882 ,  2.743 ,   72.0   ,-7.095    ,-2.137   ,    14.75  ,-0.255     ,471.263 ,   47.25  ,-420.259
14 ,     1 ,     2 ,  129 ,22612 ,0.009 ,  4 ,  9.964 ,  917.789 ,-1.945 ,  2.752 ,   72.5   ,-7.213    ,-1.989   ,     6.75  ,-0.044     ,475.903 ,   48.0   ,-441.885
 9 ,     1 ,     2 ,   99 ,22953 ,0.028 , 98 , 10.036 ,  891.777 ,-2.004 ,  2.723 ,   72.75  ,-7.313    ,-1.848   ,     8.0   ,0.156      ,472.717 ,   47.25  ,-419.06
 4 ,     1 ,     2 ,   21 ,19761 ,0.007 ,  3 , 10.098 ,  883.486 ,-2.014 ,  2.718 ,   73.0   ,-7.38     ,-1.939   ,     7.75  ,0.074      ,468.117 ,   47.0   ,-415.369
13 ,     1 ,     2 ,  123 ,22349 ,0.031 ,  5 , 10.314 ,  905.618 ,-2.007 ,  2.696 ,   74.0   ,-7.617    ,-1.849   ,     8.25  ,0.158      ,478.931 ,   47.0   ,-426.687
